
/*
* company:
* author/engineer:
* creation date:
* project name:
* target devices:
* tool versions:
*
* * DESCRIPTION:
*
* * INTERFACE:
*		[port name]		- [port description]
* * inputs:
* * outputs:
*/

import reg_file_pkg::*;

module reg_file_memory #(
    parameter                   MEMORY_TYPE = REG_FILE_MEMORY_TYPE_DUAL_PORT
) (
);

    //----------------------------------------------------------
    // INTERNAL SIGNALS
    //----------------------------------------------------------


    //----------------------------------------------------------
    // OPERATION
    //----------------------------------------------------------


    //----------------------------------------------------------
    // SUBMODULES
    //----------------------------------------------------------

endmodule

