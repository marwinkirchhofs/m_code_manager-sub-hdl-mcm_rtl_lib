`ifndef _AXI_REG_FILE_PARAM_H_
`define _AXI_REG_FILE_PARAM_H_

`define AXI_LITE_REG_FILE_NUM_REGISTERS 4
`define AXI_LITE_REG_FILE_AXI_ADDR_WIDTH 8

`endif
