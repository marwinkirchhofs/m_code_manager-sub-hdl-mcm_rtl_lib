
const reg_entry_t axi_lite_reg_map_table[REG_FILE_NUM_REGISTERS] = '{
    {8'h00, MEMORY_MAPPED, NO_TRIGGER_ON_WRITE, CLEAR_ON_READ},
    {8'h04, MEMORY_MAPPED, NO_TRIGGER_ON_WRITE, CLEAR_ON_READ},
    {8'h10, NO_MEMORY_MAPPED, TRIGGER_ON_WRITE, NO_CLEAR_ON_READ},
    {8'h14, MEMORY_MAPPED, TRIGGER_ON_WRITE, NO_CLEAR_ON_READ}
};
